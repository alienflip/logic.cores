`ifndef ADDER_MODULE
`define ADDER_MODULE

module adder (
    input data_0,
    input data_1,
    output out,
    output carry
);

    

endmodule

`endif 