`ifndef AGLX_ALM_MODULE
`define AGLX_ALM_MODULE

module aglx_alm (
    input       clk,
    input [7:0] data
);

endmodule

`endif