`ifndef ADDER_MODULE
`define ADDER_MODULE

module adder (
    input carry_in,
    input data_0,
    input data_1,
    output carry_out,
    output out
);

    

endmodule

`endif 