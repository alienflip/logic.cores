`ifndef F_ADDER_MODULE
`define F_ADDER_MODULE

module f_adder (
    input carry_in,
    input data_0,
    input data_1,
    output carry_out,
    output out
);

    

endmodule

`endif 