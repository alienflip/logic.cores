`include "counter.v"
`include "mplex2_1.v"
//...

module control();

endmodule